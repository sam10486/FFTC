`timescale 1 ns/1 ps     

module horizontal_tf_fly_row2(
    Q,

    rst_n,
    clk,
    state,
    stage_counter,
    CEN
) ;

parameter S_WIDTH   = 4 ; 
parameter P_WIDTH     = 64 ;
parameter SC_WIDTH    = 3; 

output reg [P_WIDTH-1:0] Q;
input                   rst_n           ;
input                   clk             ;
input [S_WIDTH-1:0]     state           ;
input [SC_WIDTH-1:0]    stage_counter   ; 
input                   CEN             ;

reg [P_WIDTH-1:0] horizontal_factor [0:63];
reg [3:0] cnt;
reg [5:0] horizontal_factor_idx;


always @(posedge clk or posedge rst_n) begin
    if (!rst_n) begin
        horizontal_factor[0] <= 64'h0000000000000001 ; // don't work
        horizontal_factor[1] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[2] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[3] <= 64'h32709a89ff61b351 ;
        horizontal_factor[4] <= 64'hbbdfdceff9b2d4ca ;
        horizontal_factor[5] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[6] <= 64'he9bf1a633740408f ;
        horizontal_factor[7] <= 64'h32709a89ff61b351 ;
        horizontal_factor[8] <= 64'ha0ab7e95c458c04e ;
        horizontal_factor[9] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[10] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[11] <= 64'h32709a89ff61b351 ;
        horizontal_factor[12] <= 64'h75755b87f702ae1f ;
        horizontal_factor[13] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[14] <= 64'he9bf1a633740408f ;
        horizontal_factor[15] <= 64'h32709a89ff61b351 ;
        horizontal_factor[16] <= 64'h7b83abdf412342cf ;
        horizontal_factor[17] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[18] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[19] <= 64'h32709a89ff61b351 ;
        horizontal_factor[20] <= 64'hbbdfdceff9b2d4ca ;
        horizontal_factor[21] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[22] <= 64'he9bf1a633740408f ;
        horizontal_factor[23] <= 64'h32709a89ff61b351 ;
        horizontal_factor[24] <= 64'hec140825b83b7edd ;
        horizontal_factor[25] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[26] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[27] <= 64'h32709a89ff61b351 ;
        horizontal_factor[28] <= 64'h75755b87f702ae1f ;
        horizontal_factor[29] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[30] <= 64'he9bf1a633740408f ;
        horizontal_factor[31] <= 64'h32709a89ff61b351 ;
        horizontal_factor[32] <= 64'hd3946b6a55f9087f ;
        horizontal_factor[33] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[34] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[35] <= 64'h32709a89ff61b351 ;
        horizontal_factor[36] <= 64'hbbdfdceff9b2d4ca ;
        horizontal_factor[37] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[38] <= 64'he9bf1a633740408f ;
        horizontal_factor[39] <= 64'h32709a89ff61b351 ;
        horizontal_factor[40] <= 64'ha0ab7e95c458c04e ;
        horizontal_factor[41] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[42] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[43] <= 64'h32709a89ff61b351 ;
        horizontal_factor[44] <= 64'h75755b87f702ae1f ;
        horizontal_factor[45] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[46] <= 64'he9bf1a633740408f ;
        horizontal_factor[47] <= 64'h32709a89ff61b351 ;
        horizontal_factor[48] <= 64'h9a12ec57bd327ded ;
        horizontal_factor[49] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[50] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[51] <= 64'h32709a89ff61b351 ;
        horizontal_factor[52] <= 64'hbbdfdceff9b2d4ca ;
        horizontal_factor[53] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[54] <= 64'he9bf1a633740408f ;
        horizontal_factor[55] <= 64'h32709a89ff61b351 ;
        horizontal_factor[56] <= 64'hec140825b83b7edd ;
        horizontal_factor[57] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[58] <= 64'hd8452f144f2e3d4b ;
        horizontal_factor[59] <= 64'h32709a89ff61b351 ;
        horizontal_factor[60] <= 64'h75755b87f702ae1f ;
        horizontal_factor[61] <= 64'h4a3f9ccc62d9a86a ;
        horizontal_factor[62] <= 64'he9bf1a633740408f ;
        horizontal_factor[63] <= 64'h32709a89ff61b351 ;
    end 
end


always @(posedge clk or posedge rst_n) begin
    if (!rst_n) begin
        cnt <= 4'd0;
    end else begin
        if (~CEN) begin
            if (stage_counter == 3'd0) begin
                if (cnt == 4'd15) begin
                    cnt <= 4'd0;
                end else begin
                    cnt <= cnt + 4'd1;
                end
            end
        end
    end
end

always @(posedge clk or posedge rst_n) begin
    if (!rst_n) begin
        horizontal_factor_idx <= 6'd1;
    end else begin
        if (cnt == 4'd15) begin
            horizontal_factor_idx <= horizontal_factor_idx + 6'd1;
        end else begin
            horizontal_factor_idx <= horizontal_factor_idx;
        end
    end
end

always @(posedge clk or posedge rst_n) begin
    if (!rst_n) begin
        Q <= 64'd0;
    end else begin
        if (~CEN) begin
           //if (cnt >= 4'd0 && cnt <= 4'd3) begin
                Q <= horizontal_factor[horizontal_factor_idx];
            //end else begin
            //    Q <= 64'd0;
            //end 
        end
    end
end

endmodule