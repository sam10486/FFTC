 `timescale 1 ns/1 ps                                                             
 module Ctrl_PipeReg1(DC_mode_sel_Dout,
                      BU_mode_sel_Dout,
                      Mul_sel_Dout,                                               
 				      RDC_sel_Dout,
					  DC_mode_sel_in,
        			  BU_mode_sel_in,		  
 			          Mul_sel_in,                                                 
 			          RDC_sel_in,                                                 
                      rst_n,                                                      
                      clk                                                         
                      ) ;                                                         
 
 output                  DC_mode_sel_Dout ;
 output                  BU_mode_sel_Dout ; 
 output                  Mul_sel_Dout ;                                           
 output [3:0]            RDC_sel_Dout ;                                           
 
 input                   DC_mode_sel_in;
 input                   BU_mode_sel_in;
 input                   Mul_sel_in ;                                             
 input  [3:0]            RDC_sel_in ;                                             
 input                   rst_n ;                                                  
 input                   clk ;                                                    


 reg                  DC_mode_sel_D0reg ;                                         
 reg                  DC_mode_sel_D1reg ;                                         
 reg                  DC_mode_sel_D2reg ;                                         
 reg                  DC_mode_sel_D3reg ;                                         
 reg                  DC_mode_sel_D4reg ;                                         
 reg                  DC_mode_sel_D5reg ;                                         
 reg                  DC_mode_sel_D6reg ;                                         
 reg                  DC_mode_sel_D7reg ;                                         
 reg                  DC_mode_sel_D8reg ;                                         
 reg                  DC_mode_sel_D9reg ;                                         
 reg                  DC_mode_sel_D10reg ;                                        
 reg                  DC_mode_sel_D11reg ;                                        
 reg                  DC_mode_sel_D12reg ;                                        
 reg                  DC_mode_sel_D13reg ;                                        
 reg                  DC_mode_sel_D14reg ;                                        
 reg                  DC_mode_sel_D15reg ;                                        
 reg                  DC_mode_sel_D16reg ;                                        
 reg                  DC_mode_sel_D17reg ;                                        
 reg                  DC_mode_sel_D18reg ;                                        
 reg                  DC_mode_sel_D19reg ;                                        
 reg                  DC_mode_sel_D20reg ;                                        
 reg                  DC_mode_sel_D21reg ;                                        
 reg                  DC_mode_sel_D22reg ;                                        
 reg                  DC_mode_sel_D23reg ;                                        
 reg                  DC_mode_sel_D24reg ;                                        
 reg                  DC_mode_sel_D25reg ;                                        
 reg                  DC_mode_sel_D26reg ;                                        
 reg                  DC_mode_sel_D27reg ;                                        
 reg                  DC_mode_sel_D28reg ;                                        
 reg                  DC_mode_sel_D29reg ;                                        
 reg                  DC_mode_sel_D30reg ;                                        
 reg                  DC_mode_sel_D31reg ;                                        
 reg                  DC_mode_sel_D32reg ;                                        
 reg                  DC_mode_sel_D33reg ;                                        
 reg                  DC_mode_sel_D34reg ;                                        
 reg                  DC_mode_sel_D35reg ;                                        
 reg                  DC_mode_sel_D36reg ;                                        
 reg                  DC_mode_sel_D37reg ;                                        
 reg                  DC_mode_sel_D38reg ;                                        
 reg                  DC_mode_sel_D39reg ;                                        
 reg                  DC_mode_sel_D40reg ;                                        
 reg                  DC_mode_sel_D41reg ;                                        
 reg                  DC_mode_sel_D42reg ;                                        
 reg                  DC_mode_sel_D43reg ;                                        
 reg                  DC_mode_sel_D44reg ;                                        
 reg                  DC_mode_sel_D45reg ;                                        
 reg                  DC_mode_sel_Dout  ;                     
 reg                  BU_mode_sel_D0reg ;                                         
 reg                  BU_mode_sel_D1reg ;                                         
 reg                  BU_mode_sel_D2reg ;                                         
 reg                  BU_mode_sel_D3reg ;                                         
 reg                  BU_mode_sel_D4reg ;                                         
 reg                  BU_mode_sel_D5reg ;                                         
 reg                  BU_mode_sel_D6reg ;                                         
 reg                  BU_mode_sel_D7reg ;                                         
 reg                  BU_mode_sel_D8reg ;                                         
 reg                  BU_mode_sel_D9reg ;                                         
 reg                  BU_mode_sel_D10reg ;                                        
 reg                  BU_mode_sel_D11reg ;                                        
 reg                  BU_mode_sel_D12reg ;                                        
 reg                  BU_mode_sel_D13reg ;                                        
 reg                  BU_mode_sel_D14reg ;                                        
 reg                  BU_mode_sel_D15reg ;                                        
 reg                  BU_mode_sel_D16reg ;                                        
 reg                  BU_mode_sel_D17reg ;                                        
 reg                  BU_mode_sel_D18reg ;                                        
 reg                  BU_mode_sel_D19reg ;                                        
 reg                  BU_mode_sel_D20reg ;                                        
 reg                  BU_mode_sel_D21reg ;                                        
 reg                  BU_mode_sel_D22reg ;                                        
 reg                  BU_mode_sel_D23reg ;                                        
 reg                  BU_mode_sel_D24reg ;                                        
 reg                  BU_mode_sel_D25reg ;                                        
 reg                  BU_mode_sel_D26reg ;                                        
 reg                  BU_mode_sel_D27reg ;                                        
 reg                  BU_mode_sel_D28reg ;                                        
 reg                  BU_mode_sel_D29reg ;                                        
 reg                  BU_mode_sel_D30reg ;                                        
 reg                  BU_mode_sel_D31reg ;                                        
 reg                  BU_mode_sel_D32reg ;                                        
 reg                  BU_mode_sel_D33reg ;                                        
 reg                  BU_mode_sel_D34reg ;                                        
 reg                  BU_mode_sel_D35reg ;                                        
 reg                  BU_mode_sel_D36reg ;                                        
 reg                  BU_mode_sel_D37reg ;                                        
 reg                  BU_mode_sel_D38reg ;                                        
 reg                  BU_mode_sel_D39reg ;                                        
 reg                  BU_mode_sel_D40reg ;                                        
 reg                  BU_mode_sel_D41reg ;                                        
 reg                  BU_mode_sel_D42reg ;                                        
 reg                  BU_mode_sel_D43reg ;                                        
 reg                  BU_mode_sel_D44reg ;                                        
 reg                  BU_mode_sel_D45reg ;                                        
 reg                  BU_mode_sel_Dout  ; 
 reg                  Mul_sel_D0reg ;                                             
 reg                  Mul_sel_D1reg ;                                             
 reg                  Mul_sel_D2reg ;                                             
 reg                  Mul_sel_D3reg ;                                             
 reg                  Mul_sel_D4reg ;                                             
 reg                  Mul_sel_Dout ;                                              
 reg [3:0]            RDC_sel_D0reg ;                                             
 reg [3:0]            RDC_sel_D1reg ;                                             
 reg [3:0]            RDC_sel_D2reg ;                                             
 reg [3:0]            RDC_sel_D3reg ;                                             
 reg [3:0]            RDC_sel_D4reg ;                                             
 reg [3:0]            RDC_sel_D5reg ;                                             
 reg [3:0]            RDC_sel_D6reg ;                                             
 reg [3:0]            RDC_sel_D7reg ;                                             
 reg [3:0]            RDC_sel_Dout ;                                              

 
 //mode_sel, Mul_sel delay 4 cycles and RDC_sel, FFT_FSmode_sel  delay 7 cycles   
 	always @(posedge clk or negedge rst_n) begin                                    
 		if(~rst_n) begin                                                                                                           
 			Mul_sel_D0reg <= 1'd0 ;                                                 
 			Mul_sel_D1reg <= 1'd0 ;                                                 
 			Mul_sel_D2reg <= 1'd0 ;                                                 
 			Mul_sel_D3reg <= 1'd0 ;                                                 
 			Mul_sel_D4reg <= 1'd0 ;                                                 
 			Mul_sel_Dout  <= 1'd0 ;                                                  
 			RDC_sel_D0reg <= 4'd0 ;                                                 
 			RDC_sel_D1reg <= 4'd0 ;                                                 
 			RDC_sel_D2reg <= 4'd0 ;                                                 
 			RDC_sel_D3reg <= 4'd0 ;                                                 
 			RDC_sel_D4reg <= 4'd0 ;                                                 
 			RDC_sel_D5reg <= 4'd0 ;                                                 
 			RDC_sel_D6reg <= 4'd0 ;                                                 
 			RDC_sel_D7reg <= 4'd0 ;                                                 
 			RDC_sel_Dout <= 4'd0 ;
            //			
 			DC_mode_sel_D0reg   <= 1'd0;                                            
 			DC_mode_sel_D1reg   <= 1'd0;                                            
 			DC_mode_sel_D2reg   <= 1'd0;                                            
 			DC_mode_sel_D3reg   <= 1'd0;                                            
 			DC_mode_sel_D4reg   <= 1'd0;                                            
 			DC_mode_sel_D5reg   <= 1'd0;                                            
 			DC_mode_sel_D6reg   <= 1'd0;                                            
 			DC_mode_sel_D7reg   <= 1'd0;                                            
 			DC_mode_sel_D8reg   <= 1'd0;                                            
 			DC_mode_sel_D9reg   <= 1'd0;                                            
 			DC_mode_sel_D10reg  <= 1'd0;                                            
 			DC_mode_sel_D11reg  <= 1'd0;                                            
 			DC_mode_sel_D12reg  <= 1'd0;                                            
 			DC_mode_sel_D13reg  <= 1'd0;                                            
 			DC_mode_sel_D14reg  <= 1'd0;                                            
 			DC_mode_sel_D15reg  <= 1'd0;                                            
 			DC_mode_sel_D16reg  <= 1'd0;                                            
 			DC_mode_sel_D17reg  <= 1'd0;                                            
 			DC_mode_sel_D18reg  <= 1'd0;                                            
 			DC_mode_sel_D19reg  <= 1'd0;                                            
 			DC_mode_sel_D20reg  <= 1'd0;                                            
 			DC_mode_sel_D21reg  <= 1'd0;                                            
 			DC_mode_sel_D22reg  <= 1'd0;                                            
 			DC_mode_sel_D23reg  <= 1'd0;                                            
 			DC_mode_sel_D24reg  <= 1'd0;                                            
 			DC_mode_sel_D25reg  <= 1'd0;                                            
 			DC_mode_sel_D26reg  <= 1'd0;                                            
 			DC_mode_sel_D27reg  <= 1'd0;                                            
 			DC_mode_sel_D28reg  <= 1'd0;                                            
 			DC_mode_sel_D29reg  <= 1'd0;                                            
 			DC_mode_sel_D30reg  <= 1'd0;                                            
 			DC_mode_sel_D31reg  <= 1'd0;                                            
 			DC_mode_sel_D32reg  <= 1'd0;                                            
 			DC_mode_sel_D33reg  <= 1'd0;                                            
 			DC_mode_sel_D34reg  <= 1'd0;                                            
 			DC_mode_sel_D35reg  <= 1'd0;                                            
 			DC_mode_sel_D36reg  <= 1'd0;                                            
 			DC_mode_sel_D37reg  <= 1'd0;                                            
 			DC_mode_sel_D38reg  <= 1'd0;                                            
 			DC_mode_sel_D39reg  <= 1'd0;                                            
 			DC_mode_sel_D40reg  <= 1'd0;                                            
 			DC_mode_sel_D41reg  <= 1'd0;                                            
 			DC_mode_sel_D42reg  <= 1'd0;                                            
 			DC_mode_sel_D43reg  <= 1'd0;                                            
 			DC_mode_sel_D44reg  <= 1'd0;                                            
 			DC_mode_sel_D45reg  <= 1'd0;                                            
 			DC_mode_sel_Dout    <= 1'd0;                          			
			//
 			BU_mode_sel_D0reg   <= 1'd0;                                            
 			BU_mode_sel_D1reg   <= 1'd0;                                            
 			BU_mode_sel_D2reg   <= 1'd0;                                            
 			BU_mode_sel_D3reg   <= 1'd0;                                            
 			BU_mode_sel_D4reg   <= 1'd0;                                            
 			BU_mode_sel_D5reg   <= 1'd0;                                            
 			BU_mode_sel_D6reg   <= 1'd0;                                            
 			BU_mode_sel_D7reg   <= 1'd0;                                            
 			BU_mode_sel_D8reg   <= 1'd0;                                            
 			BU_mode_sel_D9reg   <= 1'd0;                                            
 			BU_mode_sel_D10reg  <= 1'd0;                                             
 			BU_mode_sel_D11reg  <= 1'd0;                                             
 			BU_mode_sel_D12reg  <= 1'd0;                                             
 			BU_mode_sel_D13reg  <= 1'd0;                                             
 			BU_mode_sel_D14reg  <= 1'd0;                                             
 			BU_mode_sel_D15reg  <= 1'd0;                                             
 			BU_mode_sel_D16reg  <= 1'd0;                                             
 			BU_mode_sel_D17reg  <= 1'd0;                                             
 			BU_mode_sel_D18reg  <= 1'd0;                                             
 			BU_mode_sel_D19reg  <= 1'd0;                                             
 			BU_mode_sel_D20reg  <= 1'd0;                                             
 			BU_mode_sel_D21reg  <= 1'd0;                                             
 			BU_mode_sel_D22reg  <= 1'd0;                                             
 			BU_mode_sel_D23reg  <= 1'd0;                                             
 			BU_mode_sel_D24reg  <= 1'd0;                                             
 			BU_mode_sel_D25reg  <= 1'd0;                                             
 			BU_mode_sel_D26reg  <= 1'd0;                                             
 			BU_mode_sel_D27reg  <= 1'd0;                                             
 			BU_mode_sel_D28reg  <= 1'd0;                                             
 			BU_mode_sel_D29reg  <= 1'd0;                                             
 			BU_mode_sel_D30reg  <= 1'd0;                                             
 			BU_mode_sel_D31reg  <= 1'd0;                                             
 			BU_mode_sel_D32reg  <= 1'd0;                                             
 			BU_mode_sel_D33reg  <= 1'd0;                                             
 			BU_mode_sel_D34reg  <= 1'd0;                                             
 			BU_mode_sel_D35reg  <= 1'd0;                                             
 			BU_mode_sel_D36reg  <= 1'd0;                                             
 			BU_mode_sel_D37reg  <= 1'd0;                                             
 			BU_mode_sel_D38reg  <= 1'd0;                                             
 			BU_mode_sel_D39reg  <= 1'd0;                                             
 			BU_mode_sel_D40reg  <= 1'd0;                                             
 			BU_mode_sel_D41reg  <= 1'd0;                                             
 			BU_mode_sel_D42reg  <= 1'd0;                                             
 			BU_mode_sel_D43reg  <= 1'd0;                                             
 			BU_mode_sel_D44reg  <= 1'd0;                                             
 			BU_mode_sel_D45reg  <= 1'd0;                                             
 			BU_mode_sel_Dout    <= 1'd0;                                             			
 		end                                                                         
 		else begin                                                                                                                                                                        
 			Mul_sel_D0reg <= Mul_sel_in ;                                           
 			Mul_sel_D1reg <= Mul_sel_D0reg ;                                        
 			Mul_sel_D2reg <= Mul_sel_D1reg ;                                        
 			Mul_sel_D3reg <= Mul_sel_D2reg ;                                        
 			Mul_sel_D4reg <= Mul_sel_D3reg ;                                        
 			Mul_sel_Dout <= Mul_sel_D4reg ;                                         
 			//                                                                      
 			RDC_sel_D0reg <= RDC_sel_in ;                                           
 			RDC_sel_D1reg <= RDC_sel_D0reg ;                                        
 			RDC_sel_D2reg <= RDC_sel_D1reg ;                                        
 			RDC_sel_D3reg <= RDC_sel_D2reg ;                                        
 			RDC_sel_D4reg <= RDC_sel_D3reg ;                                        
 			RDC_sel_D5reg <= RDC_sel_D4reg ;                                        
 			RDC_sel_D6reg <= RDC_sel_D5reg ;                                        
 			RDC_sel_D7reg <= RDC_sel_D6reg ;                                        
 			RDC_sel_Dout <= RDC_sel_D7reg ;
			//
 			DC_mode_sel_D0reg   <= DC_mode_sel_in;                                  
 			DC_mode_sel_D1reg   <= DC_mode_sel_D0reg;                               
 			DC_mode_sel_D2reg   <= DC_mode_sel_D1reg;                               
 			DC_mode_sel_D3reg   <= DC_mode_sel_D2reg;                               
 			DC_mode_sel_D4reg   <= DC_mode_sel_D3reg;                               
 			DC_mode_sel_D5reg   <= DC_mode_sel_D4reg;                               
 			DC_mode_sel_D6reg   <= DC_mode_sel_D5reg;                               
 			DC_mode_sel_D7reg   <= DC_mode_sel_D6reg;                               
 			DC_mode_sel_D8reg   <= DC_mode_sel_D7reg;                               
 			DC_mode_sel_D9reg   <= DC_mode_sel_D8reg;                               
 			DC_mode_sel_D10reg  <= DC_mode_sel_D9reg;                               
 			DC_mode_sel_D11reg  <= DC_mode_sel_D10reg;                              
 			DC_mode_sel_D12reg  <= DC_mode_sel_D11reg;                              
 			DC_mode_sel_D13reg  <= DC_mode_sel_D12reg;                              
 			DC_mode_sel_D14reg  <= DC_mode_sel_D13reg;                              
 			DC_mode_sel_D15reg  <= DC_mode_sel_D14reg;                              
 			DC_mode_sel_D16reg  <= DC_mode_sel_D15reg;                              
 			DC_mode_sel_D17reg  <= DC_mode_sel_D16reg;                              
 			DC_mode_sel_D18reg  <= DC_mode_sel_D17reg;                              
 			DC_mode_sel_D19reg  <= DC_mode_sel_D18reg;                              
 			DC_mode_sel_D20reg  <= DC_mode_sel_D19reg;                              
 			DC_mode_sel_D21reg  <= DC_mode_sel_D20reg;                              
 			DC_mode_sel_D22reg  <= DC_mode_sel_D21reg;                              
 			DC_mode_sel_D23reg  <= DC_mode_sel_D22reg;                              
 			DC_mode_sel_D24reg  <= DC_mode_sel_D23reg;                              
 			DC_mode_sel_D25reg  <= DC_mode_sel_D24reg;                              
 			DC_mode_sel_D26reg  <= DC_mode_sel_D25reg;                              
 			DC_mode_sel_D27reg  <= DC_mode_sel_D26reg;                              
 			DC_mode_sel_D28reg  <= DC_mode_sel_D27reg;                              
 			DC_mode_sel_D29reg  <= DC_mode_sel_D28reg;                              
 			DC_mode_sel_D30reg  <= DC_mode_sel_D29reg;                              
 			DC_mode_sel_D31reg  <= DC_mode_sel_D30reg;                              
 			DC_mode_sel_D32reg  <= DC_mode_sel_D31reg;                              
 			DC_mode_sel_D33reg  <= DC_mode_sel_D32reg;                              
 			DC_mode_sel_D34reg  <= DC_mode_sel_D33reg;                              
 			DC_mode_sel_D35reg  <= DC_mode_sel_D34reg;                              
 			DC_mode_sel_D36reg  <= DC_mode_sel_D35reg;                              
 			DC_mode_sel_D37reg  <= DC_mode_sel_D36reg;                              
 			DC_mode_sel_D38reg  <= DC_mode_sel_D37reg;                              
 			DC_mode_sel_D39reg  <= DC_mode_sel_D38reg;                              
 			DC_mode_sel_D40reg  <= DC_mode_sel_D39reg;                              
 			DC_mode_sel_D41reg  <= DC_mode_sel_D40reg;                              
 			DC_mode_sel_D42reg  <= DC_mode_sel_D41reg;                              
 			DC_mode_sel_D43reg  <= DC_mode_sel_D42reg;                              
 			DC_mode_sel_D44reg  <= DC_mode_sel_D43reg;                              
 			DC_mode_sel_D45reg  <= DC_mode_sel_D44reg;                              
 			DC_mode_sel_Dout    <= DC_mode_sel_D45reg;               			
            //
 			BU_mode_sel_D0reg  <= BU_mode_sel_in;                                   
 			BU_mode_sel_D1reg  <= BU_mode_sel_D0reg;                                
 			BU_mode_sel_D2reg  <= BU_mode_sel_D1reg;                                
 			BU_mode_sel_D3reg  <= BU_mode_sel_D2reg;                                
 			BU_mode_sel_D4reg  <= BU_mode_sel_D3reg;                                
 			BU_mode_sel_D5reg  <= BU_mode_sel_D4reg;                                
 			BU_mode_sel_D6reg  <= BU_mode_sel_D5reg;                                
 			BU_mode_sel_D7reg  <= BU_mode_sel_D6reg;                                
 			BU_mode_sel_D8reg  <= BU_mode_sel_D7reg;                                
 			BU_mode_sel_D9reg  <= BU_mode_sel_D8reg;                                
 			BU_mode_sel_D10reg <= BU_mode_sel_D9reg;                                
 			BU_mode_sel_D11reg <= BU_mode_sel_D10reg;                               
 			BU_mode_sel_D12reg <= BU_mode_sel_D11reg;                               
 			BU_mode_sel_D13reg <= BU_mode_sel_D12reg;                               
 			BU_mode_sel_D14reg <= BU_mode_sel_D13reg;                               
 			BU_mode_sel_D15reg <= BU_mode_sel_D14reg;                               
 			BU_mode_sel_D16reg <= BU_mode_sel_D15reg;                               
 			BU_mode_sel_D17reg <= BU_mode_sel_D16reg;                               
 			BU_mode_sel_D18reg <= BU_mode_sel_D17reg;                               
 			BU_mode_sel_D19reg <= BU_mode_sel_D18reg;                               
 			BU_mode_sel_D20reg <= BU_mode_sel_D19reg;                               
 			BU_mode_sel_D21reg <= BU_mode_sel_D20reg;                               
 			BU_mode_sel_D22reg <= BU_mode_sel_D21reg;                               
 			BU_mode_sel_D23reg <= BU_mode_sel_D22reg;                               
 			BU_mode_sel_D24reg <= BU_mode_sel_D23reg;                               
 			BU_mode_sel_D25reg <= BU_mode_sel_D24reg;                               
 			BU_mode_sel_D26reg <= BU_mode_sel_D25reg;                               
 			BU_mode_sel_D27reg <= BU_mode_sel_D26reg;                               
 			BU_mode_sel_D28reg <= BU_mode_sel_D27reg;                               
 			BU_mode_sel_D29reg <= BU_mode_sel_D28reg;                               
 			BU_mode_sel_D30reg <= BU_mode_sel_D29reg;                               
 			BU_mode_sel_D31reg <= BU_mode_sel_D30reg;                               
 			BU_mode_sel_D32reg <= BU_mode_sel_D31reg;                               
 			BU_mode_sel_D33reg <= BU_mode_sel_D32reg;                               
 			BU_mode_sel_D34reg <= BU_mode_sel_D33reg;                               
 			BU_mode_sel_D35reg <= BU_mode_sel_D34reg;                               
 			BU_mode_sel_D36reg <= BU_mode_sel_D35reg;                               
 			BU_mode_sel_D37reg <= BU_mode_sel_D36reg;                               
 			BU_mode_sel_D38reg <= BU_mode_sel_D37reg;                               
 			BU_mode_sel_D39reg <= BU_mode_sel_D38reg;                               
 			BU_mode_sel_D40reg <= BU_mode_sel_D39reg;                               
 			BU_mode_sel_D41reg <= BU_mode_sel_D40reg;                               
 			BU_mode_sel_D42reg <= BU_mode_sel_D41reg;                               
 			BU_mode_sel_D43reg <= BU_mode_sel_D42reg;                               
 			BU_mode_sel_D44reg <= BU_mode_sel_D43reg;                               
 			BU_mode_sel_D45reg <= BU_mode_sel_D44reg;                               
 			BU_mode_sel_Dout   <= BU_mode_sel_D45reg;                               			
 		end                                                                         
 	end                                                                             
 endmodule                                                                        
