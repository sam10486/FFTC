`timescale 1 ns/1 ps                                                     
//5-th pipeline                                                          
module Radix16_Pipe(RA0_out,                                             
			        RA1_out,                                              
			        RA2_out,                                              
			        RA3_out,                                              
			        RA4_out,                                              
			        RA5_out,                                              
			        RA6_out,                                              
			        RA7_out,                                              
			        RA8_out,                                              
			        RA9_out,                                              
			        RA10_out,                                             
			        RA11_out,                                             
			        RA12_out,                                             
			        RA13_out,                                             
			        RA14_out,                                             
			        RA15_out,                                             
                    RA0_in,                                              
			        RA1_in,                                               
			        RA2_in,                                               
			        RA3_in,                                               
			        RA4_in,                                               
			        RA5_in,                                               
			        RA6_in,                                               
			        RA7_in,                                               
			        RA8_in,                                               
			        RA9_in,                                               
			        RA10_in,                                              
			        RA11_in,                                              
			        RA12_in,                                              
			        RA13_in,                                              
			        RA14_in,                                              
			        RA15_in,                                              
		            N_in,
                    BU_mode_sel,					
                    rst_n,                                               
                    clk                                                  
                    ) ;                                                  
                                                                         
parameter P_WIDTH     = 64 ;                                             
parameter D_WIDTH     = 192 ;                                            
                                                                         
output[P_WIDTH-1:0] RA0_out ;                                            
output[P_WIDTH-1:0] RA1_out ;                                            
output[P_WIDTH-1:0] RA2_out ;                                            
output[P_WIDTH-1:0] RA3_out ;                                            
output[P_WIDTH-1:0] RA4_out ;                                            
output[P_WIDTH-1:0] RA5_out ;                                            
output[P_WIDTH-1:0] RA6_out ;                                            
output[P_WIDTH-1:0] RA7_out ;                                            
output[P_WIDTH-1:0] RA8_out ;                                            
output[P_WIDTH-1:0] RA9_out ;                                            
output[P_WIDTH-1:0] RA10_out ;                                           
output[P_WIDTH-1:0] RA11_out ;                                           
output[P_WIDTH-1:0] RA12_out ;                                           
output[P_WIDTH-1:0] RA13_out ;                                           
output[P_WIDTH-1:0] RA14_out ;                                           
output[P_WIDTH-1:0] RA15_out ;                                           
                                                                         
input [P_WIDTH-1:0] RA0_in ;                                             
input [P_WIDTH-1:0] RA1_in ;                                             
input [P_WIDTH-1:0] RA2_in ;                                             
input [P_WIDTH-1:0] RA3_in ;                                             
input [P_WIDTH-1:0] RA4_in ;                                             
input [P_WIDTH-1:0] RA5_in ;                                             
input [P_WIDTH-1:0] RA6_in ;                                             
input [P_WIDTH-1:0] RA7_in ;                                             
input [P_WIDTH-1:0] RA8_in ;                                             
input [P_WIDTH-1:0] RA9_in ;                                             
input [P_WIDTH-1:0] RA10_in ;                                            
input [P_WIDTH-1:0] RA11_in ;                                            
input [P_WIDTH-1:0] RA12_in ;                                            
input [P_WIDTH-1:0] RA13_in ;                                            
input [P_WIDTH-1:0] RA14_in ;                                            
input [P_WIDTH-1:0] RA15_in ;                                            
input [P_WIDTH-1:0] N_in ;
input               BU_mode_sel ;                                               
input               rst_n ;                                              
input               clk ;                                                
                                                                         
//stage0                                                                 
wire  [D_WIDTH-1:0] BU_S0_0_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_0_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_1_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_1_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_2_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_2_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_3_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_3_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_4_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_4_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_5_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_5_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_6_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_6_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_7_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S0_7_R1_out_wire;                                 
wire  [D_WIDTH-1:0] R0_0;                                                
wire  [D_WIDTH-1:0] R1_0;                                                
wire  [D_WIDTH-1:0] R2_0;                                                
wire  [D_WIDTH-1:0] R3_0;                                                
wire  [D_WIDTH-1:0] R4_0;                                                
wire  [D_WIDTH-1:0] R5_0;                                                
wire  [D_WIDTH-1:0] R6_0;                                                
wire  [D_WIDTH-1:0] R7_0;                                                
wire  [D_WIDTH-1:0] R8_0;                                                
wire  [D_WIDTH-1:0] R9_0;                                                
wire  [D_WIDTH-1:0] R10_0;                                               
wire  [D_WIDTH-1:0] R11_0;                                               
wire  [D_WIDTH-1:0] R12_0;                                               
wire  [D_WIDTH-1:0] R13_0;                                               
wire  [D_WIDTH-1:0] R14_0;                                               
wire  [D_WIDTH-1:0] R15_0;                                               
 //---------------------                                                 
 //STAGE 1                                                               
wire  [D_WIDTH-1:0] R0_0_D;                                              
wire  [D_WIDTH-1:0] R1_0_D;                                              
wire  [D_WIDTH-1:0] R2_0_D;                                              
wire  [D_WIDTH-1:0] R3_0_D;                                              
wire  [D_WIDTH-1:0] R4_0_D;                                              
wire  [D_WIDTH-1:0] R5_0_D;                                              
wire  [D_WIDTH-1:0] R6_0_D;                                              
wire  [D_WIDTH-1:0] R7_0_D;                                              
wire  [D_WIDTH-1:0] R8_0_D;                                              
wire  [D_WIDTH-1:0] R9_0_D;                                              
wire  [D_WIDTH-1:0] R10_0_D;                                             
wire  [D_WIDTH-1:0] R11_0_D;                                             
wire  [D_WIDTH-1:0] R12_0_D;                                             
wire  [D_WIDTH-1:0] R13_0_D;                                             
wire  [D_WIDTH-1:0] R14_0_D;                                             
wire  [D_WIDTH-1:0] R15_0_D;                                             
wire  [D_WIDTH-1:0] BU_S1_0_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_0_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_1_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_1_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_2_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_2_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_3_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_3_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_4_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_4_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_5_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_5_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_6_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_6_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_7_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S1_7_R1_out_wire;                                 
wire  [D_WIDTH-1:0] R0_1;                                                
wire  [D_WIDTH-1:0] R1_1;                                                
wire  [D_WIDTH-1:0] R2_1;                                                
wire  [D_WIDTH-1:0] R3_1;                                                
wire  [D_WIDTH-1:0] R4_1;                                                
wire  [D_WIDTH-1:0] R5_1;                                                
wire  [D_WIDTH-1:0] R6_1;                                                
wire  [D_WIDTH-1:0] R7_1;                                                
wire  [D_WIDTH-1:0] R8_1;                                                
wire  [D_WIDTH-1:0] R9_1;                                                
wire  [D_WIDTH-1:0] R10_1;                                               
wire  [D_WIDTH-1:0] R11_1;                                               
wire  [D_WIDTH-1:0] R12_1;                                               
wire  [D_WIDTH-1:0] R13_1;                                               
wire  [D_WIDTH-1:0] R14_1;                                               
wire  [D_WIDTH-1:0] R15_1;                                               
 //STAGE 2                                                               
wire  [D_WIDTH-1:0] R0_1_D;                                              
wire  [D_WIDTH-1:0] R1_1_D;                                              
wire  [D_WIDTH-1:0] R2_1_D;                                              
wire  [D_WIDTH-1:0] R3_1_D;                                              
wire  [D_WIDTH-1:0] R4_1_D;                                              
wire  [D_WIDTH-1:0] R5_1_D;                                              
wire  [D_WIDTH-1:0] R6_1_D;                                              
wire  [D_WIDTH-1:0] R7_1_D;                                              
wire  [D_WIDTH-1:0] R8_1_D;                                              
wire  [D_WIDTH-1:0] R9_1_D;                                              
wire  [D_WIDTH-1:0] R10_1_D;                                             
wire  [D_WIDTH-1:0] R11_1_D;                                             
wire  [D_WIDTH-1:0] R12_1_D;                                             
wire  [D_WIDTH-1:0] R13_1_D;                                             
wire  [D_WIDTH-1:0] R14_1_D;                                             
wire  [D_WIDTH-1:0] R15_1_D;                                             
wire  [D_WIDTH-1:0] BU_S2_0_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_0_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_1_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_1_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_2_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_2_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_3_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_3_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_4_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_4_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_5_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_5_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_6_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_6_R1_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_7_R0_out_wire;                                 
wire  [D_WIDTH-1:0] BU_S2_7_R1_out_wire;                                 
wire  [D_WIDTH-1:0] R0_2;                                                
wire  [D_WIDTH-1:0] R1_2;                                                
wire  [D_WIDTH-1:0] R2_2;                                                
wire  [D_WIDTH-1:0] R3_2;                                                
wire  [D_WIDTH-1:0] R4_2;                                                
wire  [D_WIDTH-1:0] R5_2;                                                
wire  [D_WIDTH-1:0] R6_2;                                                
wire  [D_WIDTH-1:0] R7_2;                                                
wire  [D_WIDTH-1:0] R8_2;                                                
wire  [D_WIDTH-1:0] R9_2;                                                
wire  [D_WIDTH-1:0] R10_2;                                               
wire  [D_WIDTH-1:0] R11_2;                                               
wire  [D_WIDTH-1:0] R12_2;                                               
wire  [D_WIDTH-1:0] R13_2;                                               
wire  [D_WIDTH-1:0] R14_2;                                               
wire  [D_WIDTH-1:0] R15_2;                                               
 //STAGE 3                                                               
wire  [D_WIDTH-1:0] R0_2_D;                                              
wire  [D_WIDTH-1:0] R1_2_D;                                              
wire  [D_WIDTH-1:0] R2_2_D;                                              
wire  [D_WIDTH-1:0] R3_2_D;                                              
wire  [D_WIDTH-1:0] R4_2_D;                                              
wire  [D_WIDTH-1:0] R5_2_D;                                              
wire  [D_WIDTH-1:0] R6_2_D;                                              
wire  [D_WIDTH-1:0] R7_2_D;                                              
wire  [D_WIDTH-1:0] R8_2_D;                                              
wire  [D_WIDTH-1:0] R9_2_D;                                              
wire  [D_WIDTH-1:0] R10_2_D;                                             
wire  [D_WIDTH-1:0] R11_2_D;                                             
wire  [D_WIDTH-1:0] R12_2_D;                                             
wire  [D_WIDTH-1:0] R13_2_D;                                             
wire  [D_WIDTH-1:0] R14_2_D;                                             
wire  [D_WIDTH-1:0] R15_2_D;                                             
wire  [D_WIDTH-1:0] R0_3;                                                
wire  [D_WIDTH-1:0] R1_3;                                                
wire  [D_WIDTH-1:0] R2_3;                                                
wire  [D_WIDTH-1:0] R3_3;                                                
wire  [D_WIDTH-1:0] R4_3;                                                
wire  [D_WIDTH-1:0] R5_3;                                                
wire  [D_WIDTH-1:0] R6_3;                                                
wire  [D_WIDTH-1:0] R7_3;                                                
wire  [D_WIDTH-1:0] R8_3;                                                
wire  [D_WIDTH-1:0] R9_3;                                                
wire  [D_WIDTH-1:0] R10_3;                                               
wire  [D_WIDTH-1:0] R11_3;                                               
wire  [D_WIDTH-1:0] R12_3;                                               
wire  [D_WIDTH-1:0] R13_3;                                               
wire  [D_WIDTH-1:0] R14_3;                                               
wire  [D_WIDTH-1:0] R15_3;                                            	  
 //stage4                                                                
wire  [D_WIDTH-1:0] R0_3_D;                                              
wire  [D_WIDTH-1:0] R1_3_D;                                              
wire  [D_WIDTH-1:0] R2_3_D;                                              
wire  [D_WIDTH-1:0] R3_3_D;                                              
wire  [D_WIDTH-1:0] R4_3_D;                                              
wire  [D_WIDTH-1:0] R5_3_D;                                              
wire  [D_WIDTH-1:0] R6_3_D;                                              
wire  [D_WIDTH-1:0] R7_3_D;                                              
wire  [D_WIDTH-1:0] R8_3_D;                                              
wire  [D_WIDTH-1:0] R9_3_D;                                              
wire  [D_WIDTH-1:0] R10_3_D;                                             
wire  [D_WIDTH-1:0] R11_3_D;                                             
wire  [D_WIDTH-1:0] R12_3_D;                                             
wire  [D_WIDTH-1:0] R13_3_D;                                             
wire  [D_WIDTH-1:0] R14_3_D;                                             
wire  [D_WIDTH-1:0] R15_3_D;
//
 //Mod192_output                                                         
wire  [P_WIDTH-1:0] R0_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R1_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R2_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R3_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R4_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R5_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R6_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R7_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R8_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R9_Mod192_S_out;                                     
wire  [P_WIDTH-1:0] R10_Mod192_S_out;                                    
wire  [P_WIDTH-1:0] R11_Mod192_S_out;                                    
wire  [P_WIDTH-1:0] R12_Mod192_S_out;                                    
wire  [P_WIDTH-1:0] R13_Mod192_S_out;                                    
wire  [P_WIDTH-1:0] R14_Mod192_S_out;                                    
wire  [P_WIDTH-1:0] R15_Mod192_S_out;    

                                             
//stage 0                                                                
BU_S0 BU_S0_0(.R0_out(BU_S0_0_R0_out_wire),                              
              .R1_out(BU_S0_0_R1_out_wire),                              
              .R0_in(RA0_in),                                            
              .R1_in(RA8_in)                                             
              );                                                         
BU_S0 BU_S0_1(.R0_out(BU_S0_1_R0_out_wire),                              
              .R1_out(BU_S0_1_R1_out_wire),                              
              .R0_in(RA1_in),                                            
              .R1_in(RA9_in)                                             
              );                                                         
BU_S0 BU_S0_2(.R0_out(BU_S0_2_R0_out_wire),                              
              .R1_out(BU_S0_2_R1_out_wire),                              
              .R0_in(RA2_in),                                            
              .R1_in(RA10_in)                                            
              );                                                         
BU_S0 BU_S0_3(.R0_out(BU_S0_3_R0_out_wire),                              
              .R1_out(BU_S0_3_R1_out_wire),                              
              .R0_in(RA3_in),                                            
              .R1_in(RA11_in)                                            
              );                                                         
BU_S0 BU_S0_4(.R0_out(BU_S0_4_R0_out_wire),                              
              .R1_out(BU_S0_4_R1_out_wire),                              
              .R0_in(RA4_in),                                            
              .R1_in(RA12_in)                                            
              );                                                         
BU_S0 BU_S0_5(.R0_out(BU_S0_5_R0_out_wire),                              
              .R1_out(BU_S0_5_R1_out_wire),                              
              .R0_in(RA5_in),                                            
              .R1_in(RA13_in)                                            
              );                                                         
BU_S0 BU_S0_6(.R0_out(BU_S0_6_R0_out_wire),                              
              .R1_out(BU_S0_6_R1_out_wire),                              
              .R0_in(RA6_in),                                            
              .R1_in(RA14_in)                                            
              );                                                         
BU_S0 BU_S0_7(.R0_out(BU_S0_7_R0_out_wire),                              
              .R1_out(BU_S0_7_R1_out_wire),                              
              .R0_in(RA7_in),                                            
              .R1_in(RA15_in)                                            
              );                                                         
                                                                         
assign R0_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA0_in } : BU_S0_0_R0_out_wire;                                      
assign R1_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA1_in } : BU_S0_1_R0_out_wire;                                      
assign R2_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA2_in } : BU_S0_2_R0_out_wire;                                      
assign R3_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA3_in } : BU_S0_3_R0_out_wire;                                      
assign R4_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA4_in } : BU_S0_4_R0_out_wire;                                      
assign R5_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA5_in } : BU_S0_5_R0_out_wire;                                      
assign R6_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA6_in } : BU_S0_6_R0_out_wire;                                      
assign R7_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA7_in } : BU_S0_7_R0_out_wire;                                      
assign R8_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA8_in } : BU_S0_0_R1_out_wire;                                      
assign R9_0  = (BU_mode_sel == 1'b1) ? {128'd0 , RA9_in } : {BU_S0_1_R1_out_wire[179:0],BU_S0_1_R1_out_wire[191:180]};
assign R10_0 = (BU_mode_sel == 1'b1) ? {128'd0 , RA10_in} : {BU_S0_2_R1_out_wire[167:0],BU_S0_2_R1_out_wire[191:168]};
assign R11_0 = (BU_mode_sel == 1'b1) ? {128'd0 , RA11_in} : {BU_S0_3_R1_out_wire[155:0],BU_S0_3_R1_out_wire[191:156]};
assign R12_0 = (BU_mode_sel == 1'b1) ? {128'd0 , RA12_in} : {BU_S0_4_R1_out_wire[143:0],BU_S0_4_R1_out_wire[191:144]};
assign R13_0 = (BU_mode_sel == 1'b1) ? {128'd0 , RA13_in} : {BU_S0_5_R1_out_wire[131:0],BU_S0_5_R1_out_wire[191:132]};
assign R14_0 = (BU_mode_sel == 1'b1) ? {128'd0 , RA14_in} : {BU_S0_6_R1_out_wire[119:0],BU_S0_6_R1_out_wire[191:120]};
assign R15_0 = (BU_mode_sel == 1'b1) ? {128'd0 , RA15_in} : {BU_S0_7_R1_out_wire[107:0],BU_S0_7_R1_out_wire[191:108]};
                                                                         
 Pipe Pipe_STAGE_0(.R0_out(R0_0_D),                                      
                   .R1_out(R1_0_D),                                      
                   .R2_out(R2_0_D),                                      
                   .R3_out(R3_0_D),                                      
                   .R4_out(R4_0_D),                                      
                   .R5_out(R5_0_D),                                      
                   .R6_out(R6_0_D),                                      
                   .R7_out(R7_0_D),                                      
                   .R8_out(R8_0_D),                                      
                   .R9_out(R9_0_D),                                      
                   .R10_out(R10_0_D),                                    
                   .R11_out(R11_0_D),                                    
                   .R12_out(R12_0_D),                                    
                   .R13_out(R13_0_D),                                    
                   .R14_out(R14_0_D),                                    
                   .R15_out(R15_0_D),                                    
                   .R0_in(R0_0),                                         
                   .R1_in(R1_0),                                         
                   .R2_in(R2_0),                                         
                   .R3_in(R3_0),                                         
                   .R4_in(R4_0),                                         
                   .R5_in(R5_0),                                         
                   .R6_in(R6_0),                                         
                   .R7_in(R7_0),                                         
                   .R8_in(R8_0),                                         
                   .R9_in(R9_0),                                         
                   .R10_in(R10_0),                                       
                   .R11_in(R11_0),                                       
                   .R12_in(R12_0),                                       
                   .R13_in(R13_0),                                       
                   .R14_in(R14_0),                                       
                   .R15_in(R15_0),                                       
                   .clk(clk),                                            
                   .rst_n(rst_n)                                         
                   );                                                    
 BU BU_S1_0(.R0_out(BU_S1_0_R0_out_wire),                                
            .R1_out(BU_S1_0_R1_out_wire),                                
            .R0_in(R0_0_D),                                              
            .R1_in(R4_0_D)                                               
           );                                                            
                                                                         
 BU BU_S1_1(.R0_out(BU_S1_1_R0_out_wire),                                
            .R1_out(BU_S1_1_R1_out_wire),                                
            .R0_in(R1_0_D),                                              
            .R1_in(R5_0_D)                                               
           );                                                            
                                                                         
 BU BU_S1_2(.R0_out(BU_S1_2_R0_out_wire),                                
            .R1_out(BU_S1_2_R1_out_wire),                                
            .R0_in(R2_0_D),                                              
            .R1_in(R6_0_D)                                               
           );                                                            
                                                                         
 BU BU_S1_3(.R0_out(BU_S1_3_R0_out_wire),                                
            .R1_out(BU_S1_3_R1_out_wire),                                
            .R0_in(R3_0_D),                                              
            .R1_in(R7_0_D)                                               
           );                                                            
                                                                         
 BU BU_S1_4(.R0_out(BU_S1_4_R0_out_wire),                                
            .R1_out(BU_S1_4_R1_out_wire),                                
            .R0_in(R8_0_D),                                              
            .R1_in(R12_0_D)                                              
           );                                                            
                                                                         
 BU BU_S1_5(.R0_out(BU_S1_5_R0_out_wire),                                
            .R1_out(BU_S1_5_R1_out_wire),                                
            .R0_in(R9_0_D),                                              
            .R1_in(R13_0_D)                                              
           );                                                            
                                                                         
 BU BU_S1_6(.R0_out(BU_S1_6_R0_out_wire),                                
            .R1_out(BU_S1_6_R1_out_wire),                                
            .R0_in(R10_0_D),                                             
            .R1_in(R14_0_D)                                              
           );                                                            
                                                                         
 BU BU_S1_7(.R0_out(BU_S1_7_R0_out_wire),                                
            .R1_out(BU_S1_7_R1_out_wire),                                
            .R0_in(R11_0_D),                                             
            .R1_in(R15_0_D)                                              
           );                                                            
                                                                         
assign R0_1  = (BU_mode_sel == 1'b1) ? R0_0_D  : BU_S1_0_R0_out_wire;                                      
assign R1_1  = (BU_mode_sel == 1'b1) ? R1_0_D  : BU_S1_1_R0_out_wire;                                      
assign R2_1  = (BU_mode_sel == 1'b1) ? R2_0_D  : BU_S1_2_R0_out_wire;                                      
assign R3_1  = (BU_mode_sel == 1'b1) ? R3_0_D  : BU_S1_3_R0_out_wire;                                      
assign R4_1  = (BU_mode_sel == 1'b1) ? R4_0_D  : BU_S1_0_R1_out_wire;                                      
assign R5_1  = (BU_mode_sel == 1'b1) ? R5_0_D  : {BU_S1_1_R1_out_wire[167:0],BU_S1_1_R1_out_wire[191:168]};
assign R6_1  = (BU_mode_sel == 1'b1) ? R6_0_D  : {BU_S1_2_R1_out_wire[143:0],BU_S1_2_R1_out_wire[191:144]};
assign R7_1  = (BU_mode_sel == 1'b1) ? R7_0_D  : {BU_S1_3_R1_out_wire[119:0],BU_S1_3_R1_out_wire[191:120]};
assign R8_1  = (BU_mode_sel == 1'b1) ? R8_0_D  : BU_S1_4_R0_out_wire;                                      
assign R9_1  = (BU_mode_sel == 1'b1) ? R9_0_D  : BU_S1_5_R0_out_wire;                                      
assign R10_1 = (BU_mode_sel == 1'b1) ? R10_0_D : BU_S1_6_R0_out_wire;                                      
assign R11_1 = (BU_mode_sel == 1'b1) ? R11_0_D : BU_S1_7_R0_out_wire;                                      
assign R12_1 = (BU_mode_sel == 1'b1) ? R12_0_D : BU_S1_4_R1_out_wire;                                      
assign R13_1 = (BU_mode_sel == 1'b1) ? R13_0_D : {BU_S1_5_R1_out_wire[167:0],BU_S1_5_R1_out_wire[191:168]};
assign R14_1 = (BU_mode_sel == 1'b1) ? R14_0_D : {BU_S1_6_R1_out_wire[143:0],BU_S1_6_R1_out_wire[191:144]};
assign R15_1 = (BU_mode_sel == 1'b1) ? R15_0_D : {BU_S1_7_R1_out_wire[119:0],BU_S1_7_R1_out_wire[191:120]};
                                                                         
 Pipe Pipe_STAGE_1(.R0_out(R0_1_D),                                      
                   .R1_out(R1_1_D),                                      
                   .R2_out(R2_1_D),                                      
                   .R3_out(R3_1_D),                                      
                   .R4_out(R4_1_D),                                      
                   .R5_out(R5_1_D),                                      
                   .R6_out(R6_1_D),                                      
                   .R7_out(R7_1_D),                                      
                   .R8_out(R8_1_D),                                      
                   .R9_out(R9_1_D),                                      
                   .R10_out(R10_1_D),                                    
                   .R11_out(R11_1_D),                                    
                   .R12_out(R12_1_D),                                    
                   .R13_out(R13_1_D),                                    
                   .R14_out(R14_1_D),                                    
                   .R15_out(R15_1_D),                                    
                   .R0_in(R0_1),                                         
                   .R1_in(R1_1),                                         
                   .R2_in(R2_1),                                         
                   .R3_in(R3_1),                                         
                   .R4_in(R4_1),                                         
                   .R5_in(R5_1),                                         
                   .R6_in(R6_1),                                         
                   .R7_in(R7_1),                                         
                   .R8_in(R8_1),                                         
                   .R9_in(R9_1),                                         
                   .R10_in(R10_1),                                       
                   .R11_in(R11_1),                                       
                   .R12_in(R12_1),                                       
                   .R13_in(R13_1),                                       
                   .R14_in(R14_1),                                       
                   .R15_in(R15_1),                                       
                   .clk(clk),                                            
                   .rst_n(rst_n)                                         
                   );                                                    
                                                                         
                                                                         
 BU BU_S2_0(.R0_out(BU_S2_0_R0_out_wire),                                
            .R1_out(BU_S2_0_R1_out_wire),                                
            .R0_in(R0_1_D),                                              
            .R1_in(R2_1_D)                                               
           );                                                            
                                                                         
 BU BU_S2_1(.R0_out(BU_S2_1_R0_out_wire),                                
            .R1_out(BU_S2_1_R1_out_wire),                                
            .R0_in(R1_1_D),                                              
            .R1_in(R3_1_D)                                               
           );                                                            
                                                                         
 BU BU_S2_2(.R0_out(BU_S2_2_R0_out_wire),                                
            .R1_out(BU_S2_2_R1_out_wire),                                
            .R0_in(R4_1_D),                                              
            .R1_in(R6_1_D)                                               
           );                                                            
                                                                         
 BU BU_S2_3(.R0_out(BU_S2_3_R0_out_wire),                                
            .R1_out(BU_S2_3_R1_out_wire),                                
            .R0_in(R5_1_D),                                              
            .R1_in(R7_1_D)                                               
           );                                                            
                                                                         
 BU BU_S2_4(.R0_out(BU_S2_4_R0_out_wire),                                
            .R1_out(BU_S2_4_R1_out_wire),                                
            .R0_in(R8_1_D),                                              
            .R1_in(R10_1_D)                                              
           );                                                            
                                                                         
 BU BU_S2_5(.R0_out(BU_S2_5_R0_out_wire),                                
            .R1_out(BU_S2_5_R1_out_wire),                                
            .R0_in(R9_1_D),                                              
            .R1_in(R11_1_D)                                              
           );                                                            
                                                                         
 BU BU_S2_6(.R0_out(BU_S2_6_R0_out_wire),                                
            .R1_out(BU_S2_6_R1_out_wire),                                
            .R0_in(R12_1_D),                                             
            .R1_in(R14_1_D)                                              
           );                                                            
                                                                         
 BU BU_S2_7(.R0_out(BU_S2_7_R0_out_wire),                                
            .R1_out(BU_S2_7_R1_out_wire),                                
            .R0_in(R13_1_D),                                             
            .R1_in(R15_1_D)                                              
           );                                                            
                                                                         
assign R0_2  = BU_S2_0_R0_out_wire;                                      
assign R1_2  = BU_S2_1_R0_out_wire;                                      
assign R2_2  = BU_S2_0_R1_out_wire;                                      
assign R3_2  = {BU_S2_1_R1_out_wire[143:0],BU_S2_1_R1_out_wire[191:144]};
assign R4_2  = BU_S2_2_R0_out_wire;                                      
assign R5_2  = BU_S2_3_R0_out_wire;                                      
assign R6_2  = BU_S2_2_R1_out_wire;                                      
assign R7_2  = {BU_S2_3_R1_out_wire[143:0],BU_S2_3_R1_out_wire[191:144]};
assign R8_2  = BU_S2_4_R0_out_wire;                                      
assign R9_2  = BU_S2_5_R0_out_wire;                                      
assign R10_2 = BU_S2_4_R1_out_wire;                                      
assign R11_2 = {BU_S2_5_R1_out_wire[143:0],BU_S2_5_R1_out_wire[191:144]};
assign R12_2 = BU_S2_6_R0_out_wire;                                      
assign R13_2 = BU_S2_7_R0_out_wire;                                      
assign R14_2 = BU_S2_6_R1_out_wire;                                      
assign R15_2 = {BU_S2_7_R1_out_wire[143:0],BU_S2_7_R1_out_wire[191:144]};
                                             
                                             
 Pipe Pipe_STAGE_2(.R0_out(R0_2_D),          
                   .R1_out(R1_2_D),          
                   .R2_out(R2_2_D),          
                   .R3_out(R3_2_D),          
                   .R4_out(R4_2_D),          
                   .R5_out(R5_2_D),          
                   .R6_out(R6_2_D),          
                   .R7_out(R7_2_D),          
                   .R8_out(R8_2_D),          
                   .R9_out(R9_2_D),          
                   .R10_out(R10_2_D),        
                   .R11_out(R11_2_D),        
                   .R12_out(R12_2_D),        
                   .R13_out(R13_2_D),        
                   .R14_out(R14_2_D),        
                   .R15_out(R15_2_D),        
                   .R0_in(R0_2),             
                   .R1_in(R1_2),             
                   .R2_in(R2_2),             
                   .R3_in(R3_2),             
                   .R4_in(R4_2),             
                   .R5_in(R5_2),             
                   .R6_in(R6_2),             
                   .R7_in(R7_2),             
                   .R8_in(R8_2),             
                   .R9_in(R9_2),             
                   .R10_in(R10_2),           
                   .R11_in(R11_2),           
                   .R12_in(R12_2),           
                   .R13_in(R13_2),           
                   .R14_in(R14_2),           
                   .R15_in(R15_2),           
                   .clk(clk),                
                   .rst_n(rst_n)	          
                   );                        
                                             
 BU BU_S3_0(.R0_out(R0_3),                   
            .R1_out(R1_3),                   
            .R0_in(R0_2_D),                  
            .R1_in(R1_2_D)                   
           );                                
                                             
 BU BU_S3_1(.R0_out(R2_3),                   
            .R1_out(R3_3),                   
            .R0_in(R2_2_D),                  
            .R1_in(R3_2_D)                   
           );                                
                                             
 BU BU_S3_2(.R0_out(R4_3),                   
            .R1_out(R5_3),                   
            .R0_in(R4_2_D),                  
            .R1_in(R5_2_D)                   
           );                                
                                             
 BU BU_S3_3(.R0_out(R6_3),                   
            .R1_out(R7_3),                   
            .R0_in(R6_2_D),                  
            .R1_in(R7_2_D)                   
           );                                
                                             
 BU BU_S3_4(.R0_out(R8_3),                   
            .R1_out(R9_3),                   
            .R0_in(R8_2_D),                  
            .R1_in(R9_2_D)                   
           );                                
                                             
 BU BU_S3_5(.R0_out(R10_3),                  
            .R1_out(R11_3),                  
            .R0_in(R10_2_D),                 
            .R1_in(R11_2_D)                  
           );                                
                                             
 BU BU_S3_6(.R0_out(R12_3),                  
            .R1_out(R13_3),                  
            .R0_in(R12_2_D),                 
            .R1_in(R13_2_D)                  
           );                                
                                             
 BU BU_S3_7(.R0_out(R14_3),                  
            .R1_out(R15_3),                  
            .R0_in(R14_2_D),                 
            .R1_in(R15_2_D)                  
           );	                              
                                             
                                             
 Pipe Pipe_STAGE_3(.R0_out(R0_3_D),          
                   .R1_out(R1_3_D),          
                   .R2_out(R2_3_D),          
                   .R3_out(R3_3_D),          
                   .R4_out(R4_3_D),          
                   .R5_out(R5_3_D),          
                   .R6_out(R6_3_D),          
                   .R7_out(R7_3_D),          
                   .R8_out(R8_3_D),          
                   .R9_out(R9_3_D),          
                   .R10_out(R10_3_D),        
                   .R11_out(R11_3_D),        
                   .R12_out(R12_3_D),        
                   .R13_out(R13_3_D),        
                   .R14_out(R14_3_D),        
                   .R15_out(R15_3_D),        
                   .R0_in(R0_3),             
                   .R1_in(R1_3),             
                   .R2_in(R2_3),             
                   .R3_in(R3_3),             
                   .R4_in(R4_3),             
                   .R5_in(R5_3),             
                   .R6_in(R6_3),             
                   .R7_in(R7_3),             
                   .R8_in(R8_3),             
                   .R9_in(R9_3),             
                   .R10_in(R10_3),           
                   .R11_in(R11_3),           
                   .R12_in(R12_3),           
                   .R13_in(R13_3),           
                   .R14_in(R14_3),           
                   .R15_in(R15_3),           
                   .clk(clk),                
                   .rst_n(rst_n)	          
                   );  	 	              
                                             
 Mod192 R0_Mod192(.S_out(R0_Mod192_S_out),           
                  .A_in(R0_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );                         
                                             
 Mod192 R1_Mod192(.S_out(R1_Mod192_S_out),           
                  .A_in(R1_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	                      
                                             
 Mod192 R2_Mod192(.S_out(R2_Mod192_S_out),           
                  .A_in(R2_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	                      
                                             
 Mod192 R3_Mod192(.S_out(R3_Mod192_S_out),          
                  .A_in(R3_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );                         
 Mod192 R4_Mod192(.S_out(R4_Mod192_S_out),           
                  .A_in(R4_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );                         
 Mod192 R5_Mod192(.S_out(R5_Mod192_S_out),          
                  .A_in(R5_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );                         
 Mod192 R6_Mod192(.S_out(R6_Mod192_S_out),           
                  .A_in(R6_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );                         
 Mod192 R7_Mod192(.S_out(R7_Mod192_S_out),          
                  .A_in(R7_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	                      
 Mod192 R8_Mod192(.S_out(R8_Mod192_S_out),           
                  .A_in(R8_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	                      
 Mod192 R9_Mod192(.S_out(R9_Mod192_S_out),           
                  .A_in(R9_3_D),             
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	                      
 Mod192 R10_Mod192(.S_out(R10_Mod192_S_out),          
                  .A_in(R10_3_D),            
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	 	                  
 Mod192 R11_Mod192(.S_out(R11_Mod192_S_out),         
                  .A_in(R11_3_D),            
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	 	                  
 Mod192 R12_Mod192(.S_out(R12_Mod192_S_out),          
                  .A_in(R12_3_D),            
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );	 	                  
 Mod192 R13_Mod192(.S_out(R13_Mod192_S_out),         
                  .A_in(R13_3_D),            
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );		                  
 Mod192 R14_Mod192(.S_out(R14_Mod192_S_out),          
                  .A_in(R14_3_D),            
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );                         
 Mod192 R15_Mod192(.S_out(R15_Mod192_S_out),         
                  .A_in(R15_3_D),            
                  .N_in(N_in),               
                  .clk(clk),                 
                  .rst_n(rst_n)              
                  );

 assign RA0_out   = R0_Mod192_S_out;
 assign RA1_out   = ( BU_mode_sel == 1'b1) ? R2_Mod192_S_out : R8_Mod192_S_out;       
 assign RA2_out   = ( BU_mode_sel == 1'b1) ? R1_Mod192_S_out : R4_Mod192_S_out;       
 assign RA3_out   = ( BU_mode_sel == 1'b1) ? R3_Mod192_S_out : R12_Mod192_S_out;      
 assign RA4_out   = ( BU_mode_sel == 1'b1) ? R4_Mod192_S_out : R2_Mod192_S_out;       
 assign RA5_out   = ( BU_mode_sel == 1'b1) ? R6_Mod192_S_out : R10_Mod192_S_out;      
 assign RA6_out   = ( BU_mode_sel == 1'b1) ? R5_Mod192_S_out : R6_Mod192_S_out;       
 assign RA7_out   = ( BU_mode_sel == 1'b1) ? R7_Mod192_S_out : R14_Mod192_S_out;      
 assign RA8_out   = ( BU_mode_sel == 1'b1) ? R8_Mod192_S_out : R1_Mod192_S_out;
 assign RA9_out   = ( BU_mode_sel == 1'b1) ? R10_Mod192_S_out: R9_Mod192_S_out;       
 assign RA10_out  = ( BU_mode_sel == 1'b1) ? R9_Mod192_S_out : R5_Mod192_S_out;       
 assign RA11_out  = ( BU_mode_sel == 1'b1) ? R11_Mod192_S_out: R13_Mod192_S_out;      
 assign RA12_out  = ( BU_mode_sel == 1'b1) ? R12_Mod192_S_out: R3_Mod192_S_out;       
 assign RA13_out  = ( BU_mode_sel == 1'b1) ? R14_Mod192_S_out: R11_Mod192_S_out;      
 assign RA14_out  = ( BU_mode_sel == 1'b1) ? R13_Mod192_S_out: R7_Mod192_S_out;       
 assign RA15_out  =  R15_Mod192_S_out;



				  
endmodule                                    
